`ifndef defines_vh
`define defines_vh

// Arithmetic
`define ALU_ADD 4'd0
`define ALU_SUB 4'd1
// Logic
`define ALU_AND 4'd2

`endif
