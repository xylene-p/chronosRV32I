module MEMWBRegister(
//outputs
	WBData_out; 
	//controls to WB
	wb_sel_out; 
	register_write_enable_out; 

//inputs
	WBData_in; 
	clk; 
	rst; 
	en; 
	//controls to WB
	wb_sel_in; 
	register_write_enable_in; 
	); 



endmodule 