// Chronos ALU

`include "defines.vh"

module alu (
    // outputs
    output reg [31:0] alu_out;
    // inputs
    input      [31:0] op1, op2;
    input      [3:0]  alu_func;
    );



endmodule
