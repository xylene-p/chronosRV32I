module stage_IDEX(); 


endmodule 