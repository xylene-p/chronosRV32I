module EXMEMRegister(

	);

endmodule 