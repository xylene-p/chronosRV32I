`ALU_ADD 4'b0001;
`ALU_SUB 4'b0010;
